** Profile: "SCHEMATIC1-AC"  [ C:\Users\Patrick\Wuala\Electronics\EE3102\PSpice\filter take 2-schematic1-ac.sim ] 

** Creating circuit file "filter take 2-schematic1-ac.sim.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Local Libraries :
* From [PSPICE NETLIST] section of pspiceev.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 1s 0 
.PROBE 
.INC "filter take 2-SCHEMATIC1.net" 

.INC "filter take 2-SCHEMATIC1.als"


.END
